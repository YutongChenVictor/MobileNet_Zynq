`define     DATA_SIZE       8
`define     QUAN_SIZE       6
